use ieee;
use ieee;
