library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.ALL;
    
package lfsr_pkg is
  constant LFSR_W : natural := 11;  -- LFSR width
end lfsr_pkg;
